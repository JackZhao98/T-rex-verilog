module gameDelegate(
		    input wire collide,
		    output     gameover);
   
  assign gameover = collide;

endmodule // gameDelegate
